library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- This entity is a simple wrapper for the STUDENT_AREA entity,
--   providing I/Os to the board's LEDs, switches, and 
--   pushbuttons, debounced and clock-synchronised when needed.
-- It also includes a DATA_SOURCE that generates 32-bit unsigned
--   values for manipulation.

entity TOP_LEVEL is
    Generic (disp_delay : natural := 62500000);
    Port ( GCLK : in  STD_LOGIC; -- 125MHz global clock
			  -- Board buttons
           BTN : in  STD_LOGIC_VECTOR (3 downto 0);
			  -- Board switches
           SW : in  STD_LOGIC_VECTOR (1 downto 0);
			  -- Board LEDs
           LED : out  STD_LOGIC_VECTOR (3 downto 0));
end TOP_LEVEL;

architecture Behavioral of TOP_LEVEL is

signal btn_db : STD_LOGIC_VECTOR (3 downto 0); 

-- Internal control signals for the data_source component
signal rst_source, en_source : STD_LOGIC;
signal source_data : STD_LOGIC_VECTOR (31 downto 0);

--attribute keep : string;
--attribute keep of source_data : signal is "true";
--attribute keep of rst_source : signal is "true";
--attribute keep of en_source : signal is "true";


begin

-- Debouncers and synchronisers for the
--   (active high) user buttons. The outputs will be
--   active-high and synchronous to the 125MHZ clock.
debouncers: for i in 0 to 3 generate
	button_debouncer : entity work.Debouncer 
	PORT MAP(
		CLK => GCLK,
		Sig => BTN(i),
		Deb_Sig => btn_db(i) 
	);
end generate;

-- This entity will contain the work to be carried out
--   for each task. Note that some I/Os might not be needed.	
STUDENT_AREA_component: entity work.STUDENT_AREA 
GENERIC MAP (disp_delay => disp_delay)
PORT MAP(
	CLK_125MHZ => GCLK,
	USER_PB => btn_db, 		   
	SWITCHES => SW,  	   -- Not debounced
	LED_DISPLAY => LED,
	-- Control signals for the data source
	RST_SOURCE => rst_source,
	EN_SOURCE => en_source,
	SOURCE_DATA => source_data
);

-- This component will generate data for manipulation in the
--   STUDENT_AREA component. Its control signals, including
--   the clock, are generated by the STUDENT_AREA component.
-- Note that the circuit has a maximum operating frequency of
--   5MHz. The EN input can be used to put the circuit on hold. 
DATA_SOURCE_component: entity work.DATA_SOURCE 
GENERIC MAP (data_size => 16,
             num_samples => 64)
PORT MAP(
	CLK => GCLK,
	RST => rst_source,
	EN => en_source,
	DATA_OUT => source_data
);

end Behavioral;

